 
 
module system_DE2;
  reg visual_null;
 
  test_VGA  test_VGA ();
 
 
endmodule
